----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:15:55 05/09/2016 
-- Design Name: 
-- Module Name:    SEU30 - arq_SEU30 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;


entity SEU30 is
    Port ( SEU30 : in  STD_LOGIC_VECTOR (29 downto 0);
           SEU32 : out  STD_LOGIC_VECTOR (31 downto 0));
end SEU30;

architecture arq_SEU30 of SEU30 is

begin
process(SEU30)
	begin
		if(SEU30(29) = '1')then
			SEU32(29 downto 0) <= SEU30;
			SEU32(31 downto 30) <= (others=>'1');
		else
			SEU32(29 downto 0) <= SEU30;
			SEU32(31 downto 30) <= (others=>'0');
		end if;
	end process;


end arq_SEU30;

